/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : mux2to1                                                      **
 **                                                                          **
 ******************************************************************************/

module mux2to1( s,
                x,
                y,
                m);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  s;
   input  x;
   input  y;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output m;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_2;
   wire s_LOGISIM_NET_3;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_NET_0                    = x;
   assign s_LOGISIM_NET_1                    = y;
   assign s_LOGISIM_NET_2                    = s;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign m                                  = s_LOGISIM_NET_3;

   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   Multiplexer_2      MUX_1 (.Enable(1'b1),
                             .MuxIn_0(s_LOGISIM_NET_0),
                             .MuxIn_1(s_LOGISIM_NET_1),
                             .MuxOut(s_LOGISIM_NET_3),
                             .Sel(s_LOGISIM_NET_2));



endmodule
